module moduleName (
	input wire [3:0]adress,
	output reg [16:0]data
);
	[3:0]reg reg_file[0:15];
endmodule