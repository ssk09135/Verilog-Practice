module adder_8bit (
	data_1,
	data_2,
	data_out
);
	input wire [3:0]data_1;
	input wire data_2;
	output reg data_out

endmodule