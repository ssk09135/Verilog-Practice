module UART_SHIFT (
    input clk,
    input reset,
    input tx_en,
    input [7:0]tx_data
);
    always @(posedge clk posedge reset) begin
        if (reset) begin
            
        
        end
        else begin
       
        end
    end



    
endmodule